`timescale 1ns/100ps
`define CLK_PERIOD 10